-- Bouncing Ball Video 
--
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;
LIBRARY lpm;
USE lpm.lpm_components.ALL;

PACKAGE de0core IS
	COMPONENT vga_sync
 		PORT(clock_25Mhz, red, green, blue	: IN	STD_LOGIC;
         	red_out, green_out, blue_out	: OUT 	STD_LOGIC;
			horiz_sync_out, vert_sync_out	: OUT 	STD_LOGIC;
			pixel_row, pixel_column			: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
	END COMPONENT;
END de0core;

			-- Bouncing Ball Video 
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_SIGNED.all;
LIBRARY work;
USE work.de0core.all;

ENTITY ball IS
Generic(ADDR_WIDTH: integer := 12; DATA_WIDTH: integer := 1);

   PORT(SIGNAL PB1, PB2, Clock 			: IN std_logic;
        SIGNAL Red,Green,Blue 			: OUT std_logic;
        SIGNAL Horiz_sync,Vert_sync		: OUT std_logic);		
END ball;

architecture behavior of ball is

			-- Video Display Signals   
SIGNAL Red_Data, Green_Data, Blue_Data, vert_sync_int,
		reset, Ball_on, Direction			: std_logic;
SIGNAL Size 								: std_logic_vector(9 DOWNTO 0);  
SIGNAL Ball_Y_motion 						: std_logic_vector(9 DOWNTO 0);
SIGNAL Ball_Y_pos          : std_logic_vector(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(320,10);
SIGNAL Ball_X_pos				: std_logic_vector(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(220,10);
SIGNAL pixel_row, pixel_column				: std_logic_vector(9 DOWNTO 0); 

BEGIN           
   SYNC: vga_sync
 		PORT MAP(clock_25Mhz => clock, 
				red => red_data, green => green_data, blue => blue_data,	
    	     	red_out => red, green_out => green, blue_out => blue,
			 	horiz_sync_out => horiz_sync, vert_sync_out => vert_sync_int,
			 	pixel_row => pixel_row, pixel_column => pixel_column);

Size <= CONV_STD_LOGIC_VECTOR(8,10);
Ball_X_pos <= CONV_STD_LOGIC_VECTOR(320,10);

		-- need internal copy of vert_sync to read
vert_sync <= vert_sync_int;

		-- Colors for pixel data on video signal
Red_Data <=  ball_on;
		-- Turn off Green and Blue when displaying ball
Green_Data <= '0';
Blue_Data <=  '0';

RGB_Display: Process (Ball_X_pos, Ball_Y_pos, pixel_column, pixel_row, Size)
BEGIN
			-- Set Ball_on ='1' to display ball
 IF ('0' & Ball_X_pos <= pixel_column + Size) AND
 			-- compare positive numbers only
 	(Ball_X_pos + Size >= '0' & pixel_column) AND
 	('0' & Ball_Y_pos <= pixel_row + Size) AND
 	(Ball_Y_pos + Size >= '0' & pixel_row ) THEN
 		Ball_on <= '1';
 	ELSE
 		Ball_on <= '0';
END IF;
END process RGB_Display;

Move_Ball: process
VARIABLE time_something : integer range 0 to 120 := 0;
BEGIN
			-- Move ball once every vertical sync
	
	
	WAIT UNTIL vert_sync_int'event and vert_sync_int = '1';
	
		IF PB1 = '0' THEN
			time_something := 90;
		ELSIF time_something > 0 THEN
			time_something := time_something - 1;
		END IF;
		
		IF Ball_Y_pos <= Size THEN
			Ball_Y_motion <=  CONV_STD_LOGIC_VECTOR(1,10);
			
		ELSIF time_something > 85 THEN
			Ball_Y_motion <= -CONV_STD_LOGIC_VECTOR(3,10);
			
		ELSIF time_something > 80 THEN
			Ball_Y_motion <= -CONV_STD_LOGIC_VECTOR(2,10);
		
		ELSIF time_something > 75 THEN
			Ball_Y_motion <= -CONV_STD_LOGIC_VECTOR(1,10);
		
		ELSIF time_something > 70 or (('0' & Ball_Y_pos) >= CONV_STD_LOGIC_VECTOR(480,10) - Size) THEN
			Ball_Y_motion <=  CONV_STD_LOGIC_VECTOR(0,10);

		ELSIF time_something > 65 THEN
			Ball_Y_motion <=  CONV_STD_LOGIC_VECTOR(1,10);
		
		ELSIF time_something > 60 THEN
			Ball_Y_motion <=  CONV_STD_LOGIC_VECTOR(2,10);
		
		ELSIF time_something > 50 THEN
			Ball_Y_motion <=  CONV_STD_LOGIC_VECTOR(3,10);
		
		ELSIF time_something > 0 THEN
			Ball_Y_motion <=  CONV_STD_LOGIC_VECTOR(4,10);
		
		END IF;
		
		--IF PB2 = '0' THEN
			--Ball_Y_motion <= CONV_STD_LOGIC_VECTOR(2,10);
		--ELSIF PB1 = '0' THEN
--			Ball_Y_motion <= - CONV_STD_LOGIC_VECTOR(2,10);
--		ELSE
--			Ball_Y_motion <= CONV_STD_LOGIC_VECTOR(0,10);
--		END IF;
		
			-- Bounce off top or bottom of screen
			--IF ('0' & Ball_Y_pos) >= CONV_STD_LOGIC_VECTOR(480,10) - Size THEN
				--Ball_Y_motion <= - CONV_STD_LOGIC_VECTOR(2,10);
			--ELSIF Ball_Y_pos <= Size THEN
				--Ball_Y_motion <= CONV_STD_LOGIC_VECTOR(2,10);
			--END IF;
			
			-- Compute next ball Y position
				Ball_Y_pos <= Ball_Y_pos + Ball_Y_motion;
END process Move_Ball;

END behavior;

